library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.Matrixform.all;
  
entity Sbox is
	Port(
    clk               : in std_logic;
    reset              : in std_logic; 
    inputmatrix       : in  matrix ;
    outputmatrix      : out matrix 	);
end entity;

  
architecture rtl of Sbox is
       
	    signal smatrix : matrix;
 
  
begin
  
    process(clk) 
    begin
        if rising_edge(Clk) then
            if reset = '0' then
                
            else
                for i in 0 to 3 loop
					for j in 0 to 3 loop
					   case inputmatrix(i,j) is
							when x"00" => smatrix(i,j) <= x"63";
							when x"01" => smatrix(i,j) <= x"7c";
							when x"02" => smatrix(i,j) <= x"77";
							when x"03" => smatrix(i,j) <= x"7b";
							when x"04" => smatrix(i,j) <= x"f2";
							when x"05" => smatrix(i,j) <= x"6b";
							when x"06" => smatrix(i,j) <= x"6f";
							when x"07" => smatrix(i,j) <= x"c5";
							when x"08" => smatrix(i,j) <= x"30";
							when x"09" => smatrix(i,j) <= x"01";
							when x"0a" => smatrix(i,j) <= x"67";
							when x"0b" => smatrix(i,j) <= x"2b";
							when x"0c" => smatrix(i,j) <= x"fe";
							when x"0d" => smatrix(i,j) <= x"d7";
							when x"0e" => smatrix(i,j) <= x"ab";
							when x"0f" => smatrix(i,j) <= x"76";
							when x"10" => smatrix(i,j) <= x"ca";
							when x"11" => smatrix(i,j) <= x"82";
							when x"12" => smatrix(i,j) <= x"c9";
							when x"13" => smatrix(i,j) <= x"7d";
							when x"14" => smatrix(i,j) <= x"fa";
							when x"15" => smatrix(i,j) <= x"59";
							when x"16" => smatrix(i,j) <= x"47";
							when x"17" => smatrix(i,j) <= x"f0";
							when x"18" => smatrix(i,j) <= x"ad";
							when x"19" => smatrix(i,j) <= x"d4";
							when x"1a" => smatrix(i,j) <= x"a2";
							when x"1b" => smatrix(i,j) <= x"af";
							when x"1c" => smatrix(i,j) <= x"9c";
							when x"1d" => smatrix(i,j)<= x"a4";
							when x"1e" => smatrix(i,j) <= x"72";
							when x"1f" => smatrix(i,j) <= x"c0";
							when x"20" => smatrix(i,j) <= x"b7";
							when x"21" => smatrix(i,j) <= x"fd";
							when x"22" => smatrix(i,j) <= x"93";
							when x"23" => smatrix(i,j) <= x"26";
							when x"24" => smatrix(i,j) <= x"36";
							when x"25" => smatrix(i,j) <= x"3f";
							when x"26" => smatrix(i,j) <= x"f7";
							when x"27" => smatrix(i,j) <= x"cc";
							when x"28" => smatrix(i,j) <= x"34";
							when x"29" => smatrix(i,j) <= x"a5";
							when x"2a" => smatrix(i,j) <= x"e5";
							when x"2b" => smatrix(i,j) <= x"f1";
							when x"2c" => smatrix(i,j) <= x"71";
							when x"2d" => smatrix(i,j) <= x"d8";
							when x"2e" => smatrix(i,j) <= x"31";
							when x"2f" => smatrix(i,j) <= x"15";
							when x"30" => smatrix(i,j) <= x"04";
							when x"31" => smatrix(i,j) <= x"c7";
							when x"32" => smatrix(i,j) <= x"23";
							when x"33" => smatrix(i,j) <= x"c3";
							when x"34" => smatrix(i,j) <= x"18";
							when x"35" => smatrix(i,j) <= x"96";
							when x"36" => smatrix(i,j) <= x"05";
							when x"37" => smatrix(i,j) <= x"9a";
							when x"38" => smatrix(i,j) <= x"07";
							when x"39" => smatrix(i,j) <= x"12";
							when x"3a" => smatrix(i,j) <= x"80";
							when x"3b" => smatrix(i,j) <= x"e2";
							when x"3c" => smatrix(i,j) <= x"eb";
							when x"3d" => smatrix(i,j) <= x"27";
							when x"3e" => smatrix(i,j) <= x"b2";
							when x"3f" => smatrix(i,j) <= x"75";
							when x"40" => smatrix(i,j) <= x"09";
							when x"41" => smatrix(i,j) <= x"83";
							when x"42" => smatrix(i,j) <= x"2c";
							when x"43" => smatrix(i,j) <= x"1a";
							when x"44" => smatrix(i,j) <= x"1b";
							when x"45" => smatrix(i,j) <= x"6e";
							when x"46" => smatrix(i,j) <= x"5a";
							when x"47" => smatrix(i,j) <= x"a0";
							when x"48" => smatrix(i,j) <= x"52";
							when x"49" => smatrix(i,j) <= x"3b";
							when x"4a" => smatrix(i,j) <= x"d6";
							when x"4b" => smatrix(i,j) <= x"b3";
							when x"4c" => smatrix(i,j) <= x"29";
							when x"4d" => smatrix(i,j) <= x"e3";
							when x"4e" => smatrix(i,j) <= x"2f";
							when x"4f" => smatrix(i,j) <= x"84";
							when x"50" => smatrix(i,j) <= x"53";
							when x"51" => smatrix(i,j) <= x"d1";
							when x"52" => smatrix(i,j) <= x"00";
							when x"53" => smatrix(i,j) <= x"ed";
							when x"54" => smatrix(i,j) <= x"20";
							when x"55" => smatrix(i,j) <= x"fc";
							when x"56" => smatrix(i,j) <= x"b1";
							when x"57" => smatrix(i,j) <= x"5b";
							when x"58" => smatrix(i,j) <= x"6a";
							when x"59" => smatrix(i,j) <= x"cb";
							when x"5a" => smatrix(i,j) <= x"be";
							when x"5b" => smatrix(i,j) <= x"39";
							when x"5c" => smatrix(i,j) <= x"4a";
							when x"5d" => smatrix(i,j) <= x"4c";
							when x"5e" => smatrix(i,j) <= x"58";
							when x"5f" => smatrix(i,j) <= x"cf";
							when x"60" => smatrix(i,j) <= x"d0";
							when x"61" => smatrix(i,j) <= x"ef";
							when x"62" => smatrix(i,j) <= x"aa";
							when x"63" => smatrix(i,j) <= x"fb";
							when x"64" => smatrix(i,j) <= x"43";
							when x"65" => smatrix(i,j) <= x"4d";
							when x"66" => smatrix(i,j) <= x"33";
							when x"67" => smatrix(i,j) <= x"85";
							when x"68" => smatrix(i,j) <= x"45";
							when x"69" => smatrix(i,j) <= x"f9";
							when x"6a" => smatrix(i,j) <= x"02";
							when x"6b" => smatrix(i,j) <= x"7f";
							when x"6c" => smatrix(i,j) <= x"50";
							when x"6d" => smatrix(i,j) <= x"3c";
							when x"6e" => smatrix(i,j) <= x"9f";
							when x"6f" => smatrix(i,j) <= x"a8";
							when x"70" => smatrix(i,j) <= x"51";
							when x"71" => smatrix(i,j) <= x"a3";
							when x"72" => smatrix(i,j) <= x"40";
							when x"73" => smatrix(i,j) <= x"8f";
							when x"74" => smatrix(i,j) <= x"92";
							when x"75" => smatrix(i,j) <= x"9d";
							when x"76" => smatrix(i,j) <= x"38";
							when x"77" => smatrix(i,j) <= x"f5";
							when x"78" => smatrix(i,j) <= x"bc";
							when x"79" => smatrix(i,j) <= x"b6";
							when x"7a" => smatrix(i,j) <= x"da";
							when x"7b" => smatrix(i,j) <= x"21";
							when x"7c" => smatrix(i,j) <= x"10";
							when x"7d" => smatrix(i,j) <= x"ff";
							when x"7e" => smatrix(i,j) <= x"f3";
							when x"7f" => smatrix(i,j) <= x"d2";
							when x"80" => smatrix(i,j) <= x"cd";
							when x"81" => smatrix(i,j) <= x"0c";
							when x"82" => smatrix(i,j) <= x"13";
							when x"83" => smatrix(i,j) <= x"ec";
							when x"84" => smatrix(i,j) <= x"5f";
							when x"85" => smatrix(i,j) <= x"97";
							when x"86" => smatrix(i,j) <= x"44";
							when x"87" => smatrix(i,j) <= x"17";
							when x"88" => smatrix(i,j) <= x"c4";
							when x"89" => smatrix(i,j) <= x"a7";
							when x"8a" => smatrix(i,j) <= x"7e";
							when x"8b" => smatrix(i,j) <= x"3d";
							when x"8c" => smatrix(i,j) <= x"64";
							when x"8d" => smatrix(i,j) <= x"5d";
							when x"8e" => smatrix(i,j) <= x"19";
							when x"8f" => smatrix(i,j) <= x"73";
							when x"90" => smatrix(i,j) <= x"60";
							when x"91" => smatrix(i,j) <= x"81";
							when x"92" => smatrix(i,j) <= x"4f";
							when x"93" => smatrix(i,j) <= x"dc";
							when x"94" => smatrix(i,j) <= x"22";
							when x"95" => smatrix(i,j) <= x"2a";
							when x"96" => smatrix(i,j) <= x"90";
							when x"97" => smatrix(i,j) <= x"88";
							when x"98" => smatrix(i,j) <= x"46";
							when x"99" => smatrix(i,j) <= x"ee";
							when x"9a" => smatrix(i,j) <= x"b8";
							when x"9b" => smatrix(i,j) <= x"14";
							when x"9c" => smatrix(i,j) <= x"de";
							when x"9d" => smatrix(i,j) <= x"5e";
							when x"9e" => smatrix(i,j) <= x"0b";
							when x"9f" => smatrix(i,j) <= x"db";
							when x"a0" => smatrix(i,j) <= x"e0";
							when x"a1" => smatrix(i,j) <= x"32";
							when x"a2" => smatrix(i,j) <= x"3a";
							when x"a3" => smatrix(i,j) <= x"0a";
							when x"a4" => smatrix(i,j) <= x"49";
							when x"a5" => smatrix(i,j) <= x"06";
							when x"a6" => smatrix(i,j) <= x"24";
							when x"a7" => smatrix(i,j) <= x"5c";
							when x"a8" => smatrix(i,j) <= x"c2";
							when x"a9" => smatrix(i,j) <= x"d3";
							when x"aa" => smatrix(i,j) <= x"ac";
							when x"ab" => smatrix(i,j) <= x"62";
							when x"ac" => smatrix(i,j) <= x"91";
							when x"ad" => smatrix(i,j) <= x"95";
							when x"ae" => smatrix(i,j) <= x"e4";
							when x"af" => smatrix(i,j) <= x"79";
							when x"b0" => smatrix(i,j) <= x"e7";
							when x"b1" => smatrix(i,j) <= x"c8";
							when x"b2" => smatrix(i,j) <= x"37";
							when x"b3" => smatrix(i,j) <= x"6d";
							when x"b4" => smatrix(i,j) <= x"8d";
							when x"b5" => smatrix(i,j) <= x"d5";
							when x"b6" => smatrix(i,j) <= x"4e";
							when x"b7" => smatrix(i,j) <= x"a9";
							when x"b8" => smatrix(i,j) <= x"6c";
							when x"b9" => smatrix(i,j) <= x"56";
							when x"ba" => smatrix(i,j) <= x"f4";
							when x"bb" => smatrix(i,j) <= x"ea";
							when x"bc" => smatrix(i,j) <= x"65";
							when x"bd" => smatrix(i,j) <= x"7a";
							when x"be" => smatrix(i,j) <= x"ae";
							when x"bf" => smatrix(i,j) <= x"08";
							when x"c0" => smatrix(i,j) <= x"ba";
							when x"c1" => smatrix(i,j) <= x"78";
							when x"c2" => smatrix(i,j) <= x"25";
							when x"c3" => smatrix(i,j) <= x"2e";
							when x"c4" => smatrix(i,j) <= x"1c";
							when x"c5" => smatrix(i,j) <= x"a6";
							when x"c6" => smatrix(i,j) <= x"b4";
							when x"c7" => smatrix(i,j) <= x"c6";
							when x"c8" => smatrix(i,j) <= x"e8";
							when x"c9" => smatrix(i,j) <= x"dd";
							when x"ca" => smatrix(i,j) <= x"74";
							when x"cb" => smatrix(i,j) <= x"1f";
							when x"cc" => smatrix(i,j) <= x"4b";
							when x"cd" => smatrix(i,j) <= x"bd";
							when x"ce" => smatrix(i,j) <= x"8b";
							when x"cf" => smatrix(i,j) <= x"8a";
							when x"d0" => smatrix(i,j) <= x"70";
							when x"d1" => smatrix(i,j) <= x"3e";
							when x"d2" => smatrix(i,j) <= x"b5";
							when x"d3" => smatrix(i,j) <= x"66";
							when x"d4" => smatrix(i,j) <= x"48";
							when x"d5" => smatrix(i,j) <= x"03";
							when x"d6" => smatrix(i,j) <= x"f6";
							when x"d7" => smatrix(i,j) <= x"0e";
							when x"d8" => smatrix(i,j) <= x"61";
							when x"d9" => smatrix(i,j) <= x"35";
							when x"da" => smatrix(i,j) <= x"57";
							when x"db" => smatrix(i,j) <= x"b9";
							when x"dc" => smatrix(i,j) <= x"86";
							when x"dd" => smatrix(i,j) <= x"c1";
							when x"de" => smatrix(i,j) <= x"1d";
							when x"df" => smatrix(i,j) <= x"9e";
							when x"e0" => smatrix(i,j) <= x"e1";
							when x"e1" => smatrix(i,j) <= x"f8";
							when x"e2" => smatrix(i,j) <= x"98";
							when x"e3" => smatrix(i,j) <= x"11";
							when x"e4" => smatrix(i,j) <= x"69";
							when x"e5" => smatrix(i,j) <= x"d9";
							when x"e6" => smatrix(i,j) <= x"8e";
							when x"e7" => smatrix(i,j) <= x"94";
							when x"e8" => smatrix(i,j) <= x"9b";
							when x"e9" => smatrix(i,j) <= x"1e";
							when x"ea" => smatrix(i,j) <= x"87";
							when x"eb" => smatrix(i,j) <= x"e9";
							when x"ec" => smatrix(i,j) <= x"ce";
							when x"ed" => smatrix(i,j) <= x"55";
							when x"ee" => smatrix(i,j) <= x"28";
							when x"ef" => smatrix(i,j) <= x"df";
							when x"f0" => smatrix(i,j) <= x"8c";
							when x"f1" => smatrix(i,j) <= x"a1";
							when x"f2" => smatrix(i,j) <= x"89";
							when x"f3" => smatrix(i,j) <= x"0d";
							when x"f4" => smatrix(i,j) <= x"bf";
							when x"f5" => smatrix(i,j) <= x"e6";
							when x"f6" => smatrix(i,j) <= x"42";
							when x"f7" => smatrix(i,j) <= x"68";
							when x"f8" => smatrix(i,j) <= x"41";
							when x"f9" => smatrix(i,j) <= x"99";
							when x"fa" => smatrix(i,j) <= x"2d";
							when x"fb" => smatrix(i,j) <= x"0f";
							when x"fc" => smatrix(i,j) <= x"b0";
							when x"fd" => smatrix(i,j) <= x"54";
							when x"fe" => smatrix(i,j) <= x"bb";
							when x"ff" => smatrix(i,j) <= x"16";
							when others => null; 
						end case;
					end loop;
                end loop;
            end if;
        end if;
    end process;
         outputmatrix <= smatrix;
end architecture;